`define CONST_W {{16'b0000100000000000,16'b0000000000000000}, {16'b0000000000000000,16'b0000100000000000}, {16'b0000010110101000,16'b0000010110101000}, {16'b1111101001011000,16'b0000010110101000}, {16'b0000011101100100,16'b0000001100010000}, {16'b1111110011110000,16'b0000011101100100}, {16'b0000001100010000,16'b0000011101100100}, {16'b1111100010011100,16'b0000001100010000}, {16'b0000011111011001,16'b0000000110010000}, {16'b1111111001110000,16'b0000011111011001}, {16'b0000010001110010,16'b0000011010100111}, {16'b1111100101011001,16'b0000010001110010}, {16'b0000011010100111,16'b0000010001110010}, {16'b1111101110001110,16'b0000011010100111}, {16'b0000000110010000,16'b0000011111011001}, {16'b1111100000100111,16'b0000000110010000}, {16'b0000011111110110,16'b0000000011001001}, {16'b1111111100110111,16'b0000011111110110}, {16'b0000010100010011,16'b0000011000101111}, {16'b1111100111010001,16'b0000010100010011}, {16'b0000011100001110,16'b0000001111000101}, {16'b1111110000111011,16'b0000011100001110}, {16'b0000001001010011,16'b0000011110101000}, {16'b1111100001011000,16'b0000001001010011}, {16'b0000011110101000,16'b0000001001010011}, {16'b1111110110101101,16'b0000011110101000}, {16'b0000001111000101,16'b0000011100001110}, {16'b1111100011110010,16'b0000001111000101}, {16'b0000011000101111,16'b0000010100010011}, {16'b1111101011101101,16'b0000011000101111}, {16'b0000000011001001,16'b0000011111110110}, {16'b1111100000001010,16'b0000000011001001}}